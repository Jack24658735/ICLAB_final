input [9-1:0] x;
output [5-1:0] sqrt_x;

always @* begin
    case (x)
        9'd  0: sqrt_x = 0;
        9'd  1: sqrt_x = 1;
        9'd  2: sqrt_x = 1;
        9'd  3: sqrt_x = 1;
        9'd  4: sqrt_x = 2;
        9'd  5: sqrt_x = 2;
        9'd  6: sqrt_x = 2;
        9'd  7: sqrt_x = 2;
        9'd  8: sqrt_x = 2;
        9'd  9: sqrt_x = 3;
        9'd 10: sqrt_x = 3;
        9'd 11: sqrt_x = 3;
        9'd 12: sqrt_x = 3;
        9'd 13: sqrt_x = 3;
        9'd 14: sqrt_x = 3;
        9'd 15: sqrt_x = 3;
        9'd 16: sqrt_x = 4;
        9'd 17: sqrt_x = 4;
        9'd 18: sqrt_x = 4;
        9'd 19: sqrt_x = 4;
        9'd 20: sqrt_x = 4;
        9'd 21: sqrt_x = 4;
        9'd 22: sqrt_x = 4;
        9'd 23: sqrt_x = 4;
        9'd 24: sqrt_x = 4;
        9'd 25: sqrt_x = 5;
        9'd 26: sqrt_x = 5;
        9'd 27: sqrt_x = 5;
        9'd 28: sqrt_x = 5;
        9'd 29: sqrt_x = 5;
        9'd 30: sqrt_x = 5;
        9'd 31: sqrt_x = 5;
        9'd 32: sqrt_x = 5;
        9'd 33: sqrt_x = 5;
        9'd 34: sqrt_x = 5;
        9'd 35: sqrt_x = 5;
        9'd 36: sqrt_x = 6;
        9'd 37: sqrt_x = 6;
        9'd 38: sqrt_x = 6;
        9'd 39: sqrt_x = 6;
        9'd 40: sqrt_x = 6;
        9'd 41: sqrt_x = 6;
        9'd 42: sqrt_x = 6;
        9'd 43: sqrt_x = 6;
        9'd 44: sqrt_x = 6;
        9'd 45: sqrt_x = 6;
        9'd 46: sqrt_x = 6;
        9'd 47: sqrt_x = 6;
        9'd 48: sqrt_x = 6;
        9'd 49: sqrt_x = 7;
        9'd 50: sqrt_x = 7;
        9'd 51: sqrt_x = 7;
        9'd 52: sqrt_x = 7;
        9'd 53: sqrt_x = 7;
        9'd 54: sqrt_x = 7;
        9'd 55: sqrt_x = 7;
        9'd 56: sqrt_x = 7;
        9'd 57: sqrt_x = 7;
        9'd 58: sqrt_x = 7;
        9'd 59: sqrt_x = 7;
        9'd 60: sqrt_x = 7;
        9'd 61: sqrt_x = 7;
        9'd 62: sqrt_x = 7;
        9'd 63: sqrt_x = 7;
        9'd 64: sqrt_x = 8;
        9'd 65: sqrt_x = 8;
        9'd 66: sqrt_x = 8;
        9'd 67: sqrt_x = 8;
        9'd 68: sqrt_x = 8;
        9'd 69: sqrt_x = 8;
        9'd 70: sqrt_x = 8;
        9'd 71: sqrt_x = 8;
        9'd 72: sqrt_x = 8;
        9'd 73: sqrt_x = 8;
        9'd 74: sqrt_x = 8;
        9'd 75: sqrt_x = 8;
        9'd 76: sqrt_x = 8;
        9'd 77: sqrt_x = 8;
        9'd 78: sqrt_x = 8;
        9'd 79: sqrt_x = 8;
        9'd 80: sqrt_x = 8;
        9'd 81: sqrt_x = 9;
        9'd 82: sqrt_x = 9;
        9'd 83: sqrt_x = 9;
        9'd 84: sqrt_x = 9;
        9'd 85: sqrt_x = 9;
        9'd 86: sqrt_x = 9;
        9'd 87: sqrt_x = 9;
        9'd 88: sqrt_x = 9;
        9'd 89: sqrt_x = 9;
        9'd 90: sqrt_x = 9;
        9'd 91: sqrt_x = 9;
        9'd 92: sqrt_x = 9;
        9'd 93: sqrt_x = 9;
        9'd 94: sqrt_x = 9;
        9'd 95: sqrt_x = 9;
        9'd 96: sqrt_x = 9;
        9'd 97: sqrt_x = 9;
        9'd 98: sqrt_x = 9;
        9'd 99: sqrt_x = 9;
        9'd100: sqrt_x = 10;
        9'd101: sqrt_x = 10;
        9'd102: sqrt_x = 10;
        9'd103: sqrt_x = 10;
        9'd104: sqrt_x = 10;
        9'd105: sqrt_x = 10;
        9'd106: sqrt_x = 10;
        9'd107: sqrt_x = 10;
        9'd108: sqrt_x = 10;
        9'd109: sqrt_x = 10;
        9'd110: sqrt_x = 10;
        9'd111: sqrt_x = 10;
        9'd112: sqrt_x = 10;
        9'd113: sqrt_x = 10;
        9'd114: sqrt_x = 10;
        9'd115: sqrt_x = 10;
        9'd116: sqrt_x = 10;
        9'd117: sqrt_x = 10;
        9'd118: sqrt_x = 10;
        9'd119: sqrt_x = 10;
        9'd120: sqrt_x = 10;
        9'd121: sqrt_x = 11;
        9'd122: sqrt_x = 11;
        9'd123: sqrt_x = 11;
        9'd124: sqrt_x = 11;
        9'd125: sqrt_x = 11;
        9'd126: sqrt_x = 11;
        9'd127: sqrt_x = 11;
        9'd128: sqrt_x = 11;
        9'd129: sqrt_x = 11;
        9'd130: sqrt_x = 11;
        9'd131: sqrt_x = 11;
        9'd132: sqrt_x = 11;
        9'd133: sqrt_x = 11;
        9'd134: sqrt_x = 11;
        9'd135: sqrt_x = 11;
        9'd136: sqrt_x = 11;
        9'd137: sqrt_x = 11;
        9'd138: sqrt_x = 11;
        9'd139: sqrt_x = 11;
        9'd140: sqrt_x = 11;
        9'd141: sqrt_x = 11;
        9'd142: sqrt_x = 11;
        9'd143: sqrt_x = 11;
        9'd144: sqrt_x = 12;
        9'd145: sqrt_x = 12;
        9'd146: sqrt_x = 12;
        9'd147: sqrt_x = 12;
        9'd148: sqrt_x = 12;
        9'd149: sqrt_x = 12;
        9'd150: sqrt_x = 12;
        9'd151: sqrt_x = 12;
        9'd152: sqrt_x = 12;
        9'd153: sqrt_x = 12;
        9'd154: sqrt_x = 12;
        9'd155: sqrt_x = 12;
        9'd156: sqrt_x = 12;
        9'd157: sqrt_x = 12;
        9'd158: sqrt_x = 12;
        9'd159: sqrt_x = 12;
        9'd160: sqrt_x = 12;
        9'd161: sqrt_x = 12;
        9'd162: sqrt_x = 12;
        9'd163: sqrt_x = 12;
        9'd164: sqrt_x = 12;
        9'd165: sqrt_x = 12;
        9'd166: sqrt_x = 12;
        9'd167: sqrt_x = 12;
        9'd168: sqrt_x = 12;
        9'd169: sqrt_x = 13;
        9'd170: sqrt_x = 13;
        9'd171: sqrt_x = 13;
        9'd172: sqrt_x = 13;
        9'd173: sqrt_x = 13;
        9'd174: sqrt_x = 13;
        9'd175: sqrt_x = 13;
        9'd176: sqrt_x = 13;
        9'd177: sqrt_x = 13;
        9'd178: sqrt_x = 13;
        9'd179: sqrt_x = 13;
        9'd180: sqrt_x = 13;
        9'd181: sqrt_x = 13;
        9'd182: sqrt_x = 13;
        9'd183: sqrt_x = 13;
        9'd184: sqrt_x = 13;
        9'd185: sqrt_x = 13;
        9'd186: sqrt_x = 13;
        9'd187: sqrt_x = 13;
        9'd188: sqrt_x = 13;
        9'd189: sqrt_x = 13;
        9'd190: sqrt_x = 13;
        9'd191: sqrt_x = 13;
        9'd192: sqrt_x = 13;
        9'd193: sqrt_x = 13;
        9'd194: sqrt_x = 13;
        9'd195: sqrt_x = 13;
        9'd196: sqrt_x = 14;
        9'd197: sqrt_x = 14;
        9'd198: sqrt_x = 14;
        9'd199: sqrt_x = 14;
        9'd200: sqrt_x = 14;
        9'd201: sqrt_x = 14;
        9'd202: sqrt_x = 14;
        9'd203: sqrt_x = 14;
        9'd204: sqrt_x = 14;
        9'd205: sqrt_x = 14;
        9'd206: sqrt_x = 14;
        9'd207: sqrt_x = 14;
        9'd208: sqrt_x = 14;
        9'd209: sqrt_x = 14;
        9'd210: sqrt_x = 14;
        9'd211: sqrt_x = 14;
        9'd212: sqrt_x = 14;
        9'd213: sqrt_x = 14;
        9'd214: sqrt_x = 14;
        9'd215: sqrt_x = 14;
        9'd216: sqrt_x = 14;
        9'd217: sqrt_x = 14;
        9'd218: sqrt_x = 14;
        9'd219: sqrt_x = 14;
        9'd220: sqrt_x = 14;
        9'd221: sqrt_x = 14;
        9'd222: sqrt_x = 14;
        9'd223: sqrt_x = 14;
        9'd224: sqrt_x = 14;
        9'd225: sqrt_x = 15;
        9'd226: sqrt_x = 15;
        9'd227: sqrt_x = 15;
        9'd228: sqrt_x = 15;
        9'd229: sqrt_x = 15;
        9'd230: sqrt_x = 15;
        9'd231: sqrt_x = 15;
        9'd232: sqrt_x = 15;
        9'd233: sqrt_x = 15;
        9'd234: sqrt_x = 15;
        9'd235: sqrt_x = 15;
        9'd236: sqrt_x = 15;
        9'd237: sqrt_x = 15;
        9'd238: sqrt_x = 15;
        9'd239: sqrt_x = 15;
        9'd240: sqrt_x = 15;
        9'd241: sqrt_x = 15;
        9'd242: sqrt_x = 15;
        9'd243: sqrt_x = 15;
        9'd244: sqrt_x = 15;
        9'd245: sqrt_x = 15;
        9'd246: sqrt_x = 15;
        9'd247: sqrt_x = 15;
        9'd248: sqrt_x = 15;
        9'd249: sqrt_x = 15;
        9'd250: sqrt_x = 15;
        9'd251: sqrt_x = 15;
        9'd252: sqrt_x = 15;
        9'd253: sqrt_x = 15;
        9'd254: sqrt_x = 15;
        9'd255: sqrt_x = 15;
        9'd256: sqrt_x = 16;
        9'd257: sqrt_x = 16;
        9'd258: sqrt_x = 16;
        9'd259: sqrt_x = 16;
        9'd260: sqrt_x = 16;
        9'd261: sqrt_x = 16;
        9'd262: sqrt_x = 16;
        9'd263: sqrt_x = 16;
        9'd264: sqrt_x = 16;
        9'd265: sqrt_x = 16;
        9'd266: sqrt_x = 16;
        9'd267: sqrt_x = 16;
        9'd268: sqrt_x = 16;
        9'd269: sqrt_x = 16;
        9'd270: sqrt_x = 16;
        9'd271: sqrt_x = 16;
        9'd272: sqrt_x = 16;
        9'd273: sqrt_x = 16;
        9'd274: sqrt_x = 16;
        9'd275: sqrt_x = 16;
        9'd276: sqrt_x = 16;
        9'd277: sqrt_x = 16;
        9'd278: sqrt_x = 16;
        9'd279: sqrt_x = 16;
        9'd280: sqrt_x = 16;
        9'd281: sqrt_x = 16;
        9'd282: sqrt_x = 16;
        9'd283: sqrt_x = 16;
        9'd284: sqrt_x = 16;
        9'd285: sqrt_x = 16;
        9'd286: sqrt_x = 16;
        9'd287: sqrt_x = 16;
        9'd288: sqrt_x = 16;
        9'd289: sqrt_x = 17;
        9'd290: sqrt_x = 17;
        9'd291: sqrt_x = 17;
        9'd292: sqrt_x = 17;
        9'd293: sqrt_x = 17;
        9'd294: sqrt_x = 17;
        9'd295: sqrt_x = 17;
        9'd296: sqrt_x = 17;
        9'd297: sqrt_x = 17;
        9'd298: sqrt_x = 17;
        9'd299: sqrt_x = 17;
        9'd300: sqrt_x = 17;
        9'd301: sqrt_x = 17;
        9'd302: sqrt_x = 17;
        9'd303: sqrt_x = 17;
        9'd304: sqrt_x = 17;
        9'd305: sqrt_x = 17;
        9'd306: sqrt_x = 17;
        9'd307: sqrt_x = 17;
        9'd308: sqrt_x = 17;
        9'd309: sqrt_x = 17;
        9'd310: sqrt_x = 17;
        9'd311: sqrt_x = 17;
        9'd312: sqrt_x = 17;
        9'd313: sqrt_x = 17;
        9'd314: sqrt_x = 17;
        9'd315: sqrt_x = 17;
        9'd316: sqrt_x = 17;
        9'd317: sqrt_x = 17;
        9'd318: sqrt_x = 17;
        9'd319: sqrt_x = 17;
        9'd320: sqrt_x = 17;
        9'd321: sqrt_x = 17;
        9'd322: sqrt_x = 17;
        9'd323: sqrt_x = 17;
        9'd324: sqrt_x = 18;
        9'd325: sqrt_x = 18;
        9'd326: sqrt_x = 18;
        9'd327: sqrt_x = 18;
        9'd328: sqrt_x = 18;
        9'd329: sqrt_x = 18;
        9'd330: sqrt_x = 18;
        9'd331: sqrt_x = 18;
        9'd332: sqrt_x = 18;
        9'd333: sqrt_x = 18;
        9'd334: sqrt_x = 18;
        9'd335: sqrt_x = 18;
        9'd336: sqrt_x = 18;
        9'd337: sqrt_x = 18;
        9'd338: sqrt_x = 18;
        9'd339: sqrt_x = 18;
        9'd340: sqrt_x = 18;
        9'd341: sqrt_x = 18;
        9'd342: sqrt_x = 18;
        9'd343: sqrt_x = 18;
        9'd344: sqrt_x = 18;
        9'd345: sqrt_x = 18;
        9'd346: sqrt_x = 18;
        9'd347: sqrt_x = 18;
        9'd348: sqrt_x = 18;
        9'd349: sqrt_x = 18;
        9'd350: sqrt_x = 18;
        9'd351: sqrt_x = 18;
        9'd352: sqrt_x = 18;
        9'd353: sqrt_x = 18;
        9'd354: sqrt_x = 18;
        9'd355: sqrt_x = 18;
        9'd356: sqrt_x = 18;
        9'd357: sqrt_x = 18;
        9'd358: sqrt_x = 18;
        9'd359: sqrt_x = 18;
        9'd360: sqrt_x = 18;
        9'd361: sqrt_x = 19;
        9'd362: sqrt_x = 19;
        9'd363: sqrt_x = 19;
        9'd364: sqrt_x = 19;
        9'd365: sqrt_x = 19;
        9'd366: sqrt_x = 19;
        9'd367: sqrt_x = 19;
        9'd368: sqrt_x = 19;
        9'd369: sqrt_x = 19;
        9'd370: sqrt_x = 19;
        9'd371: sqrt_x = 19;
        9'd372: sqrt_x = 19;
        9'd373: sqrt_x = 19;
        9'd374: sqrt_x = 19;
        9'd375: sqrt_x = 19;
        9'd376: sqrt_x = 19;
        9'd377: sqrt_x = 19;
        9'd378: sqrt_x = 19;
        9'd379: sqrt_x = 19;
        9'd380: sqrt_x = 19;
        9'd381: sqrt_x = 19;
        9'd382: sqrt_x = 19;
        9'd383: sqrt_x = 19;
        9'd384: sqrt_x = 19;
        9'd385: sqrt_x = 19;
        9'd386: sqrt_x = 19;
        9'd387: sqrt_x = 19;
        9'd388: sqrt_x = 19;
        9'd389: sqrt_x = 19;
        9'd390: sqrt_x = 19;
        9'd391: sqrt_x = 19;
        9'd392: sqrt_x = 19;
        9'd393: sqrt_x = 19;
        9'd394: sqrt_x = 19;
        9'd395: sqrt_x = 19;
        9'd396: sqrt_x = 19;
        9'd397: sqrt_x = 19;
        9'd398: sqrt_x = 19;
        9'd399: sqrt_x = 19;
        9'd400: sqrt_x = 20;
        9'd401: sqrt_x = 20;
        9'd402: sqrt_x = 20;
        9'd403: sqrt_x = 20;
        9'd404: sqrt_x = 20;
        9'd405: sqrt_x = 20;
        9'd406: sqrt_x = 20;
        9'd407: sqrt_x = 20;
        9'd408: sqrt_x = 20;
        9'd409: sqrt_x = 20;
        9'd410: sqrt_x = 20;
        9'd411: sqrt_x = 20;
        9'd412: sqrt_x = 20;
        9'd413: sqrt_x = 20;
        9'd414: sqrt_x = 20;
        9'd415: sqrt_x = 20;
        9'd416: sqrt_x = 20;
        9'd417: sqrt_x = 20;
        9'd418: sqrt_x = 20;
        9'd419: sqrt_x = 20;
        9'd420: sqrt_x = 20;
        9'd421: sqrt_x = 20;
        9'd422: sqrt_x = 20;
        9'd423: sqrt_x = 20;
        9'd424: sqrt_x = 20;
        9'd425: sqrt_x = 20;
        9'd426: sqrt_x = 20;
        9'd427: sqrt_x = 20;
        9'd428: sqrt_x = 20;
        9'd429: sqrt_x = 20;
        9'd430: sqrt_x = 20;
        9'd431: sqrt_x = 20;
        9'd432: sqrt_x = 20;
        9'd433: sqrt_x = 20;
        9'd434: sqrt_x = 20;
        9'd435: sqrt_x = 20;
        9'd436: sqrt_x = 20;
        9'd437: sqrt_x = 20;
        9'd438: sqrt_x = 20;
        9'd439: sqrt_x = 20;
        9'd440: sqrt_x = 20;
        9'd441: sqrt_x = 21;
        9'd442: sqrt_x = 21;
        9'd443: sqrt_x = 21;
        9'd444: sqrt_x = 21;
        9'd445: sqrt_x = 21;
        9'd446: sqrt_x = 21;
        9'd447: sqrt_x = 21;
        9'd448: sqrt_x = 21;
        9'd449: sqrt_x = 21;
        9'd450: sqrt_x = 21;
        9'd451: sqrt_x = 21;
        9'd452: sqrt_x = 21;
        9'd453: sqrt_x = 21;
        9'd454: sqrt_x = 21;
        9'd455: sqrt_x = 21;
        9'd456: sqrt_x = 21;
        9'd457: sqrt_x = 21;
        9'd458: sqrt_x = 21;
        9'd459: sqrt_x = 21;
        9'd460: sqrt_x = 21;
        9'd461: sqrt_x = 21;
        9'd462: sqrt_x = 21;
        9'd463: sqrt_x = 21;
        9'd464: sqrt_x = 21;
        9'd465: sqrt_x = 21;
        9'd466: sqrt_x = 21;
        9'd467: sqrt_x = 21;
        9'd468: sqrt_x = 21;
        9'd469: sqrt_x = 21;
        9'd470: sqrt_x = 21;
        9'd471: sqrt_x = 21;
        9'd472: sqrt_x = 21;
        9'd473: sqrt_x = 21;
        9'd474: sqrt_x = 21;
        9'd475: sqrt_x = 21;
        9'd476: sqrt_x = 21;
        9'd477: sqrt_x = 21;
        9'd478: sqrt_x = 21;
        9'd479: sqrt_x = 21;
        9'd480: sqrt_x = 21;
        9'd481: sqrt_x = 21;
        9'd482: sqrt_x = 21;
        9'd483: sqrt_x = 21;
        9'd484: sqrt_x = 22;
        9'd485: sqrt_x = 22;
        9'd486: sqrt_x = 22;
        9'd487: sqrt_x = 22;
        9'd488: sqrt_x = 22;
        9'd489: sqrt_x = 22;
        9'd490: sqrt_x = 22;
        9'd491: sqrt_x = 22;
        9'd492: sqrt_x = 22;
        9'd493: sqrt_x = 22;
        9'd494: sqrt_x = 22;
        9'd495: sqrt_x = 22;
        9'd496: sqrt_x = 22;
        9'd497: sqrt_x = 22;
        9'd498: sqrt_x = 22;
        9'd499: sqrt_x = 22;
        9'd500: sqrt_x = 22;
        9'd501: sqrt_x = 22;
        9'd502: sqrt_x = 22;
        9'd503: sqrt_x = 22;
        9'd504: sqrt_x = 22;
        9'd505: sqrt_x = 22;
        9'd506: sqrt_x = 22;
        9'd507: sqrt_x = 22;
        9'd508: sqrt_x = 22;
        9'd509: sqrt_x = 22;
        9'd510: sqrt_x = 22;
        9'd511: sqrt_x = 22;
        9'd512: sqrt_x = 22;
        default: sqrt_x = 0;
    endcase
end

endmodule