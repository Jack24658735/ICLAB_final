`timescale 1ns/100ps

module test_top;

localparam END_CYCLES = 10000; // you can enlarge the cycle count limit for longer simulation
real CYCLE = 10;


endmodule