module top(
    input clk, 
    input rst_n, 
    input [8*9-1:0] pixel_in,
    output valid,
    input [8*9-1:0] pixel_out
)

endmodule